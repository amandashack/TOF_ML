* C:\Users\proxi\Downloads\MRCO_NM_Base_LTspice.asc-20231205T203243Z-001\MRCO_NM_Base_LTspice.asc
R1 N004 N001 3.08Meg
R2 N005 N004 2.43Meg
R3 N006 N005 1.75Meg
R4 N007 N006 1.25Meg
R5 N008 N007 0.897Meg
R6 N009 N008 0.664Meg
R7 N010 N009 0.528Meg
R8 N011 N010 0.446Meg
R9 N012 N011 0.457Meg
R10 N013 N012 0.483Meg
R11 N014 N013 0.528Meg
R12 N015 N014 0.577Meg
R13 N016 N015 0.621Meg
R14 N017 N016 0.650Meg
R15 N018 N017 0.657Meg
R16 N019 N018 0.639Meg
R17 N020 N019 0.593Meg
R18 N021 N020 0.520Meg
R19 N022 N021 0.422Meg
R20 N023 N022 0.305Meg
R21 N024 N023 0.178Meg
R22 N002 N024 0.048Meg
R23 N025 N002 0.072Meg
R24 N026 N025 0.167Meg
R25 N003 N026 0.220Meg
V22 0 N002 88.752
V25 0 N003 86.46000000000001
R26 N027 N003 2.13Meg
V1 0 N027 100.0
V0 0 N001 -10
* Blade 01
* Blade 02
* Blade 03
* Blade 04
* Blade 05
* Blade 06
* Blade 07
* Blade 08
* Blade 09
* Blade 10
* Blade 11
* Blade 12
* Blade 13
* Blade 14
* Blade 15
* Blade 16
* Blade 17
* Blade 18
* Blade 19
* Blade 20
* Blade 21
* Blade 22
* Blade 23
* Blade 24
* Blade 25
.op
* For NM, V22 = abs(0.11248 * abs(RetardationVal) - abs(RetardationVal))\n              V25 = abs(0.1354 * abs(RetardationVal) - abs(RetardationVal))
.backanno
.end
